module inv (
	input IN,
	output OUT );

	assign OUT = !IN;

endmodule
