`ifndef stimuli_IF
`define stimuli_IF

//`timescale 1ns / 1ps
// Not using this interface, instead connecting directly to bs_if
interface stimuli_if();

// insert signals

endinterface


`endif
